module GetKPlus(K, KPlus); 

input [1:64] K;
output [0:55] KPlus;
wire [0:55] KPlus;

assign KPlus [0:55] = {
			K[57], K[49], K[41], K[33], K[25], K[17], K[9], K[1], 
			K[58], K[50], K[42], K[34], K[26], K[18], K[10], K[2], 
			K[59], K[51], K[43], K[35], K[27], K[19], K[11], K[3], 
			K[60], K[52], K[44], K[36], K[63], K[55], K[47], K[39], 
			K[31], K[23], K[15], K[7], K[62], K[54], K[46], K[38], 
			K[30], K[22], K[14], K[6], K[61], K[53], K[45], K[37], 
			K[29], K[21], K[13], K[5], K[28], K[20], K[12], K[4]
			};
	
endmodule 