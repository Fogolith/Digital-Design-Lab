module Split_48_6(KE, Split); 
input [47:0] KE; 
output [7:0] Split [1:8]; 
wire [7:0] Split [1:8]; 

assign Split = KE; 

endmodule 